library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
	port(
		i_address : in std_logic_vector(7 downto 0);
		i_CLK     : in std_logic;
		o_instruction : out std_logic_vector(31 downto 0));
end ROM;

architecture arch_1 of ROM is

type w_array is array(0 to 28) of std_logic_vector(31 downto 0);

signal w_inst : w_array := (0 => "00100000000010000000000000000000",

 1  => "00000000000000000000000000000000",
 2  => "00000000000000000000000000000000",
 3  => "00000000000000000000000000000000",
 
 4  => "00100000000010010000000000000001",
 
 5  => "00000000000000000000000000000000",
 6  => "00000000000000000000000000000000",
 7  => "00000000000000000000000000000000",
 
 8  => "00100000000010100000000000000010",
 
 9  => "00000000000000000000000000000000",
 10 => "00000000000000000000000000000000",
 11 => "00000000000000000000000000000000",
 
 12 => "00100000000010110000000000000011",
 
 13 => "00000000000000000000000000000000",
 14 => "00000000000000000000000000000000",
 15 => "00000000000000000000000000000000",
 
 
 16 => "00100000000011000000000000000100",
 
 17 => "00000000000000000000000000000000",
 18 => "00000000000000000000000000000000",
 19 => "00000000000000000000000000000000",
 
 20 => "00010001011011000000000000011100",
 
 21 => "00000000000000000000000000000000",
 22 => "00000000000000000000000000000000",
 23 => "00000000000000000000000000000000",
 
 24 => "00000001001010100100000000100000",
 
 25 => "00000000000000000000000000000000",
 26 => "00000000000000000000000000000000",
 27 => "00000000000000000000000000000000",
 
 28 => "00000001000010110100000000100010"
 );
 
 --$zero = 00000
 --$s0 = 01000
 --$s1 = 01001
 --$s2 = 01010
 --$s3 = 01011
 --$s4 = 01100
 
begin
process (i_CLK, i_address)
begin
	if (rising_edge(i_CLK)) then
			o_instruction <= w_inst(to_integer(unsigned(i_address)));
	end if;
end process;
end arch_1;
